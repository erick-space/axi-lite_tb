

//`include "axi_lite_if.sv"
//`include "axi_stream_if.sv"


package axi_lite_pkg;



typedef enum {READ, WRITE} axi_lite_cmd_t;


endpackage // axi4lite_pkg